--===========================================================================--
--
--  S Y N T H E Z I A B L E    SWTBUG ROM   C O R E
--
--  www.OpenCores.Org - December 2002
--  This core adheres to the GNU public license  
--
-- File name      : swtbug.vhd
--
-- entity name    : rombios_rom
--
-- Purpose        : Implements a 4K x 8 ROM containing the
--                  Pyldin 601 rombios program
--                  
-- Dependencies   : ieee.Std_Logic_1164
--                  ieee.std_logic_unsigned
--                  ieee.std_logic_arith
--
-- Author         : John E. Kent      
--
--===========================================================================----
--
-- Revision History:
--
-- Date:          Revision         Author
-- 22 Sep 2002    0.1              John Kent
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rombios_rom is
port (
	addr   	: in  std_logic_vector(11 downto 0);
	data		: out std_logic_vector(7 downto 0)
);
end;

architecture basic of rombios_rom is
constant width   : integer := 8;
constant memsize : integer := 4096;

type rom_array is array(0 to memsize-1) of std_logic_vector(width-1 downto 0);

constant rom_data : rom_array := (
x"3f", x"30", x"39", x"7e", x"fa", x"02", x"0f", x"ce", x"00", x"00", x"ff", x"e6", x"2a", x"ce", x"00", x"7f", 
x"ff", x"e6", x"28", x"ce", x"37", x"37", x"ff", x"e6", x"2a", x"86", x"01", x"b7", x"e6", x"29", x"5f", x"ce", 
x"ff", x"73", x"a6", x"00", x"f7", x"e6", x"00", x"b7", x"e6", x"01", x"08", x"5c", x"c1", x"10", x"26", x"f2", 
x"ce", x"ed", x"80", x"6f", x"00", x"08", x"8c", x"f0", x"00", x"26", x"f8", x"c6", x"70", x"8e", x"fe", x"eb", 
x"ce", x"ee", x"00", x"32", x"a7", x"00", x"08", x"5a", x"26", x"f9", x"ce", x"a5", x"5a", x"bc", x"ed", x"00", 
x"27", x"1f", x"ff", x"ed", x"00", x"ce", x"01", x"00", x"6f", x"00", x"08", x"8c", x"bd", x"80", x"26", x"f8", 
x"ce", x"00", x"00", x"df", x"18", x"df", x"1a", x"ce", x"01", x"01", x"df", x"1c", x"ce", x"07", x"c5", x"df", 
x"1e", x"7f", x"e6", x"f0", x"7f", x"00", x"00", x"7f", x"00", x"01", x"7f", x"ed", x"02", x"7f", x"e6", x"c0", 
x"7c", x"e6", x"c0", x"ce", x"ff", x"6b", x"ff", x"ed", x"22", x"ee", x"02", x"ff", x"ed", x"1d", x"7f", x"ed", 
x"30", x"7f", x"ed", x"06", x"ce", x"00", x"00", x"ff", x"ee", x"14", x"ce", x"ff", x"5c", x"ff", x"ed", x"26", 
x"ce", x"bf", x"f0", x"ff", x"ed", x"0c", x"ff", x"ed", x"0e", x"86", x"60", x"b7", x"ed", x"1f", x"ce", x"ff", 
x"8a", x"ff", x"ed", x"24", x"ce", x"be", x"00", x"35", x"4f", x"5f", x"3f", x"12", x"ce", x"ff", x"d8", x"3f", 
x"23", x"c6", x"08", x"f7", x"e6", x"f0", x"ce", x"a5", x"5a", x"c5", x"04", x"27", x"03", x"ce", x"5a", x"a5", 
x"bc", x"c0", x"00", x"26", x"2b", x"ce", x"c0", x"00", x"4f", x"ab", x"00", x"08", x"8c", x"e0", x"00", x"26", 
x"f8", x"4d", x"26", x"1c", x"37", x"ce", x"c0", x"10", x"df", x"20", x"a6", x"00", x"27", x"0e", x"f6", x"e6", 
x"f0", x"ee", x"01", x"3f", x"2f", x"de", x"20", x"08", x"08", x"08", x"20", x"ec", x"bd", x"c0", x"0a", x"33", 
x"5c", x"c1", x"10", x"25", x"be", x"7f", x"e6", x"f0", x"ce", x"f0", x"00", x"4f", x"ab", x"00", x"08", x"26", 
x"fb", x"4d", x"27", x"02", x"3f", x"00", x"c6", x"02", x"3f", x"26", x"c6", x"04", x"86", x"26", x"3f", x"27", 
x"0e", x"b6", x"e6", x"d0", x"84", x"c0", x"81", x"80", x"26", x"19", x"86", x"80", x"3f", x"17", x"ce", x"ff", 
x"65", x"86", x"01", x"3f", x"17", x"4d", x"26", x"0b", x"fe", x"02", x"fe", x"8c", x"a5", x"5a", x"26", x"03", 
x"bd", x"01", x"50", x"3f", x"01", x"20", x"fc", x"f6", x"ed", x"81", x"54", x"54", x"54", x"54", x"fe", x"ee", 
x"04", x"20", x"1f", x"f6", x"ed", x"84", x"fe", x"ee", x"12", x"7d", x"e6", x"2a", x"2b", x"14", x"f6", x"ed", 
x"81", x"fe", x"ee", x"06", x"7d", x"e6", x"2b", x"2a", x"09", x"7d", x"e6", x"29", x"f6", x"ed", x"82", x"fe", 
x"ee", x"0a", x"b6", x"e6", x"f0", x"36", x"c4", x"0f", x"27", x"03", x"f7", x"e6", x"f0", x"8c", x"00", x"00", 
x"27", x"02", x"ad", x"00", x"32", x"b7", x"e6", x"f0", x"3b", x"0f", x"7c", x"00", x"00", x"30", x"ae", x"05", 
x"34", x"32", x"31", x"af", x"05", x"35", x"36", x"8d", x"3c", x"32", x"f6", x"e6", x"f0", x"37", x"16", x"54", 
x"d7", x"03", x"c6", x"ed", x"d7", x"02", x"de", x"02", x"e6", x"80", x"25", x"04", x"54", x"54", x"54", x"54", 
x"c4", x"0f", x"27", x"03", x"f7", x"e6", x"f0", x"c6", x"77", x"48", x"59", x"97", x"03", x"d7", x"02", x"de", 
x"02", x"a6", x"01", x"e6", x"00", x"27", x"02", x"8d", x"35", x"0f", x"33", x"f7", x"e6", x"f0", x"30", x"8d", 
x"04", x"7a", x"00", x"00", x"3b", x"a6", x"01", x"d6", x"05", x"97", x"05", x"e7", x"01", x"a6", x"02", x"d6", 
x"06", x"97", x"06", x"e7", x"02", x"a6", x"03", x"d6", x"07", x"97", x"07", x"e7", x"03", x"a6", x"04", x"d6", 
x"08", x"97", x"08", x"e7", x"04", x"a6", x"00", x"d6", x"04", x"97", x"04", x"e7", x"00", x"39", x"36", x"37", 
x"96", x"04", x"06", x"de", x"07", x"d6", x"05", x"96", x"06", x"0e", x"39", x"b6", x"e6", x"2a", x"88", x"08", 
x"b7", x"e6", x"2a", x"09", x"26", x"fd", x"20", x"f3", x"ce", x"00", x"00", x"bc", x"ed", x"04", x"27", x"12", 
x"c6", x"0c", x"b6", x"ed", x"04", x"bd", x"f4", x"7e", x"5c", x"b6", x"ed", x"05", x"bd", x"f4", x"7e", x"ff", 
x"ed", x"04", x"96", x"18", x"4c", x"4c", x"81", x"64", x"25", x"01", x"4f", x"97", x"18", x"26", x"48", x"3f", 
x"06", x"96", x"19", x"4c", x"81", x"3c", x"25", x"01", x"4f", x"97", x"19", x"4d", x"26", x"39", x"96", x"1a", 
x"4c", x"81", x"3c", x"25", x"01", x"4f", x"97", x"1a", x"26", x"2d", x"96", x"1b", x"4c", x"81", x"18", x"25", 
x"01", x"4f", x"97", x"1b", x"26", x"21", x"96", x"1c", x"4c", x"81", x"20", x"25", x"02", x"86", x"01", x"97", 
x"1c", x"81", x"01", x"26", x"12", x"96", x"1d", x"4c", x"81", x"0d", x"25", x"02", x"86", x"01", x"97", x"1d", 
x"81", x"01", x"26", x"03", x"7c", x"00", x"1e", x"86", x"ff", x"3f", x"17", x"7d", x"ed", x"09", x"27", x"03", 
x"7a", x"ed", x"09", x"7d", x"ed", x"0a", x"27", x"03", x"7a", x"ed", x"0a", x"7d", x"ed", x"0b", x"27", x"0a", 
x"7a", x"ed", x"0b", x"26", x"05", x"86", x"ff", x"b7", x"ed", x"31", x"39", x"7d", x"ed", x"09", x"27", x"04", 
x"b6", x"e6", x"28", x"39", x"5f", x"b6", x"e6", x"28", x"5a", x"27", x"f8", x"81", x"ff", x"27", x"f6", x"c6", 
x"1e", x"b1", x"ed", x"31", x"26", x"07", x"7d", x"ed", x"0a", x"26", x"77", x"c6", x"03", x"f7", x"ed", x"0a", 
x"b7", x"ed", x"31", x"fe", x"ed", x"0c", x"81", x"fe", x"27", x"04", x"81", x"fd", x"26", x"03", x"ff", x"ed", 
x"0e", x"08", x"8c", x"c0", x"00", x"26", x"03", x"ce", x"bf", x"f0", x"ff", x"ed", x"50", x"bc", x"ed", x"0e", 
x"27", x"50", x"f6", x"e6", x"2a", x"c5", x"08", x"27", x"1a", x"81", x"c0", x"24", x"16", x"81", x"41", x"25", 
x"12", x"81", x"5a", x"23", x"0c", x"81", x"61", x"25", x"0a", x"81", x"7a", x"23", x"04", x"81", x"80", x"25", 
x"02", x"88", x"20", x"81", x"fc", x"26", x"07", x"c8", x"08", x"f7", x"e6", x"2a", x"20", x"22", x"81", x"fb", 
x"26", x"13", x"b6", x"e6", x"29", x"88", x"01", x"b7", x"e6", x"29", x"c6", x"60", x"44", x"25", x"01", x"5f", 
x"f7", x"ed", x"1f", x"20", x"0b", x"fe", x"ed", x"0c", x"a7", x"00", x"fe", x"ed", x"50", x"ff", x"ed", x"0c", 
x"8d", x"0b", x"c6", x"03", x"f7", x"ed", x"09", x"c6", x"05", x"f7", x"ed", x"0b", x"39", x"86", x"0f", x"f6", 
x"e6", x"2b", x"c8", x"08", x"f7", x"e6", x"2b", x"f6", x"ed", x"0a", x"5a", x"01", x"26", x"fc", x"f6", x"e6", 
x"2b", x"c8", x"08", x"f7", x"e6", x"2b", x"f6", x"ed", x"0a", x"5c", x"c1", x"3c", x"26", x"fb", x"4a", x"26", 
x"de", x"39", x"0f", x"86", x"ff", x"fe", x"ed", x"0e", x"bc", x"ed", x"0c", x"27", x"02", x"a6", x"00", x"97", 
x"06", x"39", x"20", x"05", x"b1", x"ed", x"1f", x"27", x"12", x"b6", x"ed", x"1f", x"36", x"ba", x"ed", x"1d", 
x"c6", x"0a", x"8d", x"2e", x"5c", x"b6", x"ed", x"1e", x"8d", x"28", x"32", x"0e", x"01", x"0f", x"fe", x"ed", 
x"0e", x"bc", x"ed", x"0c", x"27", x"de", x"a6", x"00", x"08", x"8c", x"c0", x"00", x"26", x"03", x"ce", x"bf", 
x"f0", x"ff", x"ed", x"0e", x"97", x"06", x"fe", x"ed", x"22", x"c6", x"0a", x"a6", x"06", x"8d", x"03", x"5c", 
x"a6", x"07", x"7e", x"f4", x"7e", x"0f", x"84", x"7f", x"81", x"05", x"25", x"01", x"39", x"84", x"03", x"7f", 
x"ed", x"56", x"ff", x"ed", x"13", x"ff", x"ed", x"19", x"b7", x"ed", x"12", x"97", x"0d", x"81", x"02", x"26", 
x"0a", x"f7", x"ed", x"1b", x"c4", x"03", x"58", x"58", x"58", x"20", x"0a", x"4d", x"26", x"06", x"5d", x"27", 
x"03", x"f7", x"ed", x"1c", x"5f", x"86", x"ff", x"97", x"0c", x"de", x"0c", x"ea", x"85", x"b6", x"e6", x"29", 
x"84", x"c1", x"b7", x"e6", x"29", x"fa", x"e6", x"29", x"f7", x"e6", x"29", x"ce", x"ff", x"73", x"a6", x"06", 
x"f6", x"ed", x"12", x"c4", x"03", x"26", x"32", x"b7", x"ed", x"17", x"4c", x"4c", x"8d", x"5e", x"a6", x"01", 
x"b7", x"ed", x"18", x"4c", x"4c", x"8d", x"52", x"ee", x"10", x"ff", x"ed", x"15", x"c6", x"f0", x"f7", x"ed", 
x"13", x"86", x"00", x"b7", x"ed", x"14", x"7d", x"00", x"06", x"2a", x"06", x"f6", x"ed", x"19", x"b6", x"ed", 
x"1a", x"f7", x"ed", x"19", x"b7", x"ed", x"1a", x"20", x"12", x"8d", x"31", x"a6", x"01", x"8d", x"2a", x"f6", 
x"ed", x"13", x"b6", x"ed", x"14", x"54", x"46", x"54", x"46", x"54", x"46", x"37", x"c6", x"0d", x"8d", x"1e", 
x"5a", x"32", x"8d", x"1a", x"7d", x"00", x"06", x"2b", x"0f", x"ce", x"bf", x"a0", x"c6", x"50", x"6f", x"00", 
x"08", x"5a", x"26", x"fa", x"86", x"0c", x"3f", x"22", x"39", x"c6", x"01", x"8c", x"c6", x"06", x"f7", x"e6", 
x"00", x"b7", x"e6", x"01", x"39", x"0f", x"fe", x"ed", x"13", x"f6", x"ed", x"1b", x"b6", x"ed", x"12", x"85", 
x"03", x"26", x"03", x"f6", x"ed", x"1c", x"7e", x"ff", x"f0", x"0f", x"fe", x"ed", x"19", x"b6", x"ed", x"10", 
x"f6", x"ed", x"11", x"7e", x"ff", x"f0", x"0f", x"f1", x"ed", x"17", x"24", x"0b", x"f7", x"ed", x"11", x"b1", 
x"ed", x"18", x"24", x"03", x"b7", x"ed", x"10", x"7e", x"fa", x"bf", x"0f", x"f7", x"ed", x"1c", x"39", x"0f", 
x"7f", x"ed", x"6d", x"81", x"ff", x"27", x"56", x"81", x"80", x"27", x"65", x"4d", x"26", x"03", x"7e", x"f5", 
x"87", x"e6", x"00", x"53", x"c4", x"01", x"f7", x"ed", x"67", x"e6", x"01", x"f7", x"ed", x"68", x"e6", x"02", 
x"c4", x"01", x"f7", x"ed", x"69", x"58", x"58", x"fa", x"ed", x"67", x"f7", x"ed", x"6e", x"e6", x"03", x"f7", 
x"ed", x"6a", x"ee", x"04", x"ff", x"ed", x"6b", x"b7", x"ed", x"7b", x"84", x"7f", x"c6", x"52", x"ce", x"f6", 
x"76", x"4a", x"27", x"36", x"c6", x"57", x"ce", x"f6", x"ef", x"4a", x"27", x"2e", x"c6", x"53", x"ce", x"f5", 
x"b5", x"4a", x"27", x"26", x"c6", x"46", x"ce", x"f7", x"89", x"4a", x"27", x"1e", x"39", x"7d", x"ed", x"62", 
x"27", x"0d", x"7a", x"ed", x"62", x"26", x"08", x"b6", x"e6", x"c0", x"84", x"07", x"b7", x"e6", x"c0", x"39", 
x"7f", x"ed", x"62", x"86", x"ff", x"b7", x"ed", x"64", x"20", x"4d", x"df", x"0c", x"fe", x"ed", x"20", x"e7", 
x"51", x"de", x"0c", x"f6", x"ed", x"62", x"7f", x"ed", x"62", x"86", x"01", x"48", x"ba", x"ed", x"67", x"48", 
x"0d", x"49", x"b7", x"e6", x"c0", x"8a", x"02", x"b7", x"ed", x"63", x"b6", x"ed", x"67", x"b1", x"ed", x"64", 
x"26", x"03", x"5d", x"26", x"08", x"c6", x"00", x"4a", x"26", x"fd", x"5a", x"26", x"fa", x"ad", x"00", x"fe", 
x"ed", x"20", x"6f", x"51", x"b6", x"ed", x"67", x"b7", x"ed", x"64", x"fe", x"ed", x"26", x"a6", x"08", x"b7", 
x"ed", x"62", x"7d", x"ed", x"6d", x"27", x"02", x"8d", x"0c", x"b6", x"ed", x"6d", x"97", x"06", x"96", x"18", 
x"8b", x"0a", x"97", x"18", x"39", x"7f", x"e6", x"c0", x"86", x"01", x"b7", x"e6", x"c0", x"86", x"ff", x"b7", 
x"ed", x"61", x"86", x"03", x"b7", x"ed", x"6f", x"fe", x"ed", x"26", x"ee", x"00", x"ff", x"ed", x"70", x"c6", 
x"03", x"bd", x"f8", x"77", x"39", x"8d", x"0e", x"7d", x"ed", x"6d", x"26", x"08", x"bd", x"f6", x"dd", x"f6", 
x"ed", x"72", x"d7", x"05", x"39", x"5f", x"b6", x"ed", x"67", x"0d", x"59", x"4a", x"2a", x"fc", x"f5", x"ed", 
x"61", x"27", x"1a", x"f8", x"ed", x"61", x"f7", x"ed", x"61", x"86", x"07", x"b7", x"ed", x"6f", x"b6", x"ed", 
x"67", x"b7", x"ed", x"70", x"c6", x"02", x"bd", x"f8", x"77", x"86", x"50", x"8d", x"34", x"86", x"0f", x"b7", 
x"ed", x"6f", x"b6", x"ed", x"6e", x"b7", x"ed", x"70", x"b6", x"ed", x"68", x"7d", x"ed", x"7b", x"2a", x"01", 
x"48", x"b7", x"ed", x"71", x"c6", x"03", x"bd", x"f8", x"77", x"f6", x"ed", x"68", x"b6", x"ed", x"65", x"7d", 
x"ed", x"67", x"27", x"03", x"b6", x"ed", x"66", x"7d", x"ed", x"7b", x"2a", x"01", x"58", x"10", x"2a", x"01", 
x"40", x"4c", x"fe", x"ed", x"26", x"e6", x"00", x"53", x"54", x"54", x"54", x"54", x"5c", x"f7", x"ed", x"78", 
x"fe", x"ed", x"78", x"01", x"09", x"26", x"fc", x"4a", x"26", x"f6", x"86", x"08", x"b7", x"ed", x"6f", x"c6", 
x"01", x"bd", x"f8", x"77", x"c6", x"02", x"bd", x"f8", x"9c", x"7d", x"ed", x"6d", x"26", x"27", x"b6", x"ed", 
x"70", x"7d", x"ed", x"67", x"26", x"05", x"b7", x"ed", x"65", x"20", x"03", x"b7", x"ed", x"66", x"b6", x"ed", 
x"6f", x"84", x"60", x"81", x"60", x"26", x"0e", x"86", x"20", x"ba", x"ed", x"6d", x"b7", x"ed", x"6d", x"b6", 
x"ed", x"63", x"b7", x"e6", x"c0", x"39", x"bd", x"f5", x"c5", x"7d", x"ed", x"6d", x"27", x"01", x"39", x"86", 
x"66", x"bd", x"f8", x"43", x"fe", x"ed", x"6b", x"b6", x"e6", x"d0", x"2b", x"27", x"7f", x"ed", x"78", x"b6", 
x"e6", x"d0", x"2b", x"1f", x"7c", x"ed", x"79", x"26", x"f6", x"7c", x"ed", x"78", x"26", x"f1", x"84", x"20", 
x"27", x"2d", x"86", x"40", x"bd", x"f6", x"69", x"20", x"26", x"b6", x"e6", x"d0", x"2b", x"05", x"b6", x"e6", 
x"d0", x"2a", x"eb", x"b6", x"e6", x"d1", x"a7", x"00", x"08", x"5a", x"26", x"ed", x"b6", x"e6", x"d0", x"2b", 
x"05", x"b6", x"e6", x"d0", x"2a", x"d8", x"b6", x"e6", x"d1", x"a7", x"00", x"08", x"5a", x"26", x"ed", x"b6", 
x"ed", x"63", x"b7", x"e6", x"c0", x"c6", x"07", x"bd", x"f8", x"9c", x"7e", x"f8", x"d5", x"86", x"4a", x"b7", 
x"ed", x"6f", x"b6", x"ed", x"6e", x"b7", x"ed", x"70", x"c6", x"02", x"bd", x"f8", x"77", x"20", x"e6", x"86", 
x"05", x"b7", x"ed", x"7a", x"7a", x"ed", x"7a", x"2a", x"01", x"39", x"bd", x"f5", x"8e", x"7f", x"ed", x"6d", 
x"bd", x"f8", x"21", x"bd", x"f5", x"c5", x"7d", x"ed", x"6d", x"26", x"ee", x"8d", x"d0", x"7d", x"ed", x"6d", 
x"26", x"e7", x"86", x"45", x"bd", x"f8", x"43", x"fe", x"ed", x"6b", x"b6", x"e6", x"d0", x"2b", x"2c", x"7f", 
x"ed", x"78", x"b6", x"e6", x"d0", x"2b", x"24", x"7c", x"ed", x"79", x"26", x"f6", x"7c", x"ed", x"78", x"26", 
x"f1", x"84", x"20", x"27", x"37", x"86", x"40", x"bd", x"f6", x"69", x"20", x"30", x"b6", x"e6", x"d0", x"2b", 
x"0a", x"b6", x"e6", x"d0", x"2b", x"05", x"b6", x"e6", x"d0", x"2a", x"e6", x"a6", x"00", x"b7", x"e6", x"d1", 
x"08", x"5a", x"26", x"e8", x"b6", x"e6", x"d0", x"2b", x"0a", x"b6", x"e6", x"d0", x"2b", x"05", x"b6", x"e6", 
x"d0", x"2a", x"ce", x"a6", x"00", x"b7", x"e6", x"d1", x"08", x"5a", x"26", x"e8", x"b6", x"ed", x"63", x"b7", 
x"e6", x"c0", x"c6", x"07", x"bd", x"f8", x"9c", x"bd", x"f8", x"d5", x"b6", x"ed", x"6d", x"81", x"40", x"27", 
x"05", x"81", x"02", x"27", x"01", x"39", x"7e", x"f6", x"f4", x"86", x"05", x"b7", x"ed", x"7a", x"7a", x"ed", 
x"7a", x"2a", x"01", x"39", x"bd", x"f5", x"8e", x"7f", x"ed", x"6d", x"bd", x"f8", x"21", x"bd", x"f5", x"c5", 
x"7d", x"ed", x"6d", x"26", x"ee", x"86", x"4d", x"b7", x"ed", x"6f", x"b6", x"ed", x"6e", x"b7", x"ed", x"70", 
x"fe", x"ed", x"26", x"a6", x"02", x"b7", x"ed", x"71", x"a6", x"03", x"b7", x"ed", x"72", x"a6", x"06", x"b7", 
x"ed", x"73", x"a6", x"07", x"b7", x"ed", x"74", x"c6", x"06", x"bd", x"f8", x"77", x"fe", x"ed", x"6b", x"f6", 
x"ed", x"6a", x"58", x"58", x"b6", x"e6", x"d0", x"2b", x"22", x"b6", x"e6", x"d0", x"2b", x"1d", x"7f", x"ed", 
x"78", x"b6", x"e6", x"d0", x"2b", x"15", x"7c", x"ed", x"79", x"26", x"f6", x"7c", x"ed", x"78", x"26", x"f1", 
x"84", x"20", x"27", x"10", x"86", x"40", x"bd", x"f6", x"69", x"20", x"09", x"a6", x"00", x"b7", x"e6", x"d1", 
x"08", x"5a", x"26", x"d0", x"b6", x"ed", x"63", x"b7", x"e6", x"c0", x"c6", x"07", x"bd", x"f8", x"9c", x"bd", 
x"f8", x"d5", x"b6", x"ed", x"6d", x"81", x"40", x"27", x"05", x"81", x"02", x"27", x"01", x"39", x"7e", x"f7", 
x"8e", x"86", x"04", x"b7", x"ed", x"6f", x"b6", x"ed", x"6e", x"b7", x"ed", x"70", x"c6", x"02", x"bd", x"f8", 
x"77", x"c6", x"01", x"bd", x"f8", x"9c", x"b6", x"ed", x"6f", x"84", x"40", x"26", x"01", x"39", x"86", x"01", 
x"7e", x"f6", x"69", x"b7", x"ed", x"6f", x"b6", x"ed", x"6e", x"b7", x"ed", x"70", x"b6", x"ed", x"68", x"b7", 
x"ed", x"71", x"b6", x"ed", x"69", x"b7", x"ed", x"72", x"b6", x"ed", x"6a", x"b7", x"ed", x"73", x"fe", x"ed", 
x"26", x"a6", x"02", x"b7", x"ed", x"74", x"a6", x"03", x"b7", x"ed", x"75", x"a6", x"04", x"b7", x"ed", x"76", 
x"a6", x"05", x"b7", x"ed", x"77", x"c6", x"09", x"ce", x"ed", x"6f", x"7f", x"ed", x"78", x"b6", x"e6", x"d0", 
x"84", x"c0", x"81", x"80", x"27", x"0c", x"7a", x"ed", x"78", x"26", x"f2", x"31", x"31", x"86", x"40", x"7e", 
x"f6", x"69", x"a6", x"00", x"b7", x"e6", x"d1", x"08", x"5a", x"26", x"df", x"39", x"ce", x"ed", x"6f", x"b6", 
x"e6", x"d0", x"84", x"c0", x"81", x"c0", x"27", x"1b", x"7f", x"ed", x"78", x"b6", x"e6", x"d0", x"84", x"c0", 
x"81", x"c0", x"27", x"0f", x"7a", x"ed", x"79", x"26", x"f2", x"7a", x"ed", x"78", x"26", x"ed", x"86", x"40", 
x"7e", x"f6", x"69", x"b6", x"e6", x"d1", x"a7", x"00", x"08", x"5a", x"26", x"d3", x"b6", x"ed", x"63", x"88", 
x"02", x"b7", x"e6", x"c0", x"39", x"7d", x"ed", x"6d", x"26", x"36", x"b6", x"ed", x"6f", x"84", x"c0", x"27", 
x"2f", x"c6", x"80", x"81", x"40", x"26", x"21", x"b6", x"ed", x"70", x"c6", x"08", x"48", x"8d", x"19", x"c6", 
x"04", x"48", x"48", x"8d", x"13", x"c6", x"02", x"48", x"8d", x"0e", x"c6", x"08", x"48", x"48", x"8d", x"08", 
x"c6", x"01", x"48", x"8d", x"03", x"c6", x"10", x"48", x"24", x"06", x"fa", x"ed", x"6d", x"f7", x"ed", x"6d", 
x"39", x"37", x"8d", x"1c", x"f6", x"e6", x"29", x"58", x"24", x"03", x"73", x"ed", x"7c", x"33", x"39", x"8d", 
x"1b", x"e6", x"00", x"54", x"8d", x"0f", x"e6", x"01", x"8d", x"e7", x"46", x"5a", x"26", x"fa", x"8d", x"e1", 
x"e6", x"00", x"8c", x"c6", x"14", x"5a", x"26", x"fd", x"f6", x"ed", x"7c", x"39", x"fe", x"ed", x"24", x"f6", 
x"e6", x"29", x"2b", x"f8", x"e6", x"02", x"f7", x"ed", x"7c", x"39", x"0f", x"7c", x"00", x"18", x"8d", x"cf", 
x"0d", x"26", x"01", x"0c", x"97", x"06", x"07", x"97", x"04", x"39", x"0f", x"7c", x"00", x"18", x"8d", x"dc", 
x"0c", x"8d", x"0f", x"e6", x"01", x"44", x"8d", x"0a", x"5a", x"26", x"fa", x"53", x"fb", x"ed", x"7c", x"8d", 
x"01", x"0d", x"37", x"f6", x"e6", x"29", x"c4", x"bf", x"24", x"05", x"ca", x"40", x"73", x"ed", x"7c", x"f7", 
x"e6", x"29", x"8d", x"ac", x"33", x"39", x"7d", x"ed", x"06", x"26", x"2a", x"3f", x"11", x"81", x"fe", x"27", 
x"07", x"fe", x"ed", x"22", x"a1", x"01", x"26", x"04", x"3f", x"04", x"20", x"ef", x"fe", x"ee", x"14", x"27", 
x"22", x"e6", x"00", x"c1", x"ff", x"27", x"1c", x"11", x"27", x"08", x"08", x"e6", x"00", x"26", x"fb", x"08", 
x"20", x"ef", x"ff", x"ed", x"07", x"fe", x"ed", x"07", x"08", x"ff", x"ed", x"07", x"a6", x"00", x"b7", x"ed", 
x"06", x"27", x"c3", x"7e", x"ff", x"f4", x"b6", x"ed", x"18", x"b0", x"ed", x"10", x"4a", x"11", x"24", x"01", 
x"16", x"f7", x"ed", x"7d", x"5f", x"3f", x"20", x"81", x"c0", x"27", x"22", x"22", x"f8", x"81", x"7f", x"26", 
x"07", x"5d", x"27", x"f1", x"09", x"5a", x"20", x"11", x"f1", x"ed", x"7d", x"26", x"04", x"86", x"07", x"20", 
x"08", x"a7", x"00", x"08", x"5c", x"81", x"20", x"25", x"dc", x"3f", x"22", x"20", x"d8", x"6f", x"00", x"d7", 
x"06", x"39", x"36", x"37", x"16", x"07", x"36", x"17", x"0f", x"ff", x"ed", x"5f", x"8d", x"08", x"fe", x"ed", 
x"5f", x"32", x"06", x"33", x"32", x"39", x"0f", x"f6", x"ed", x"12", x"c4", x"03", x"26", x"21", x"7d", x"ed", 
x"56", x"27", x"43", x"fe", x"ed", x"57", x"a7", x"00", x"08", x"ff", x"ed", x"57", x"7a", x"ed", x"56", x"26", 
x"5b", x"ce", x"ed", x"59", x"e6", x"00", x"c1", x"1f", x"26", x"06", x"a6", x"01", x"b7", x"ed", x"1c", x"39", 
x"c1", x"1b", x"26", x"04", x"a6", x"01", x"20", x"29", x"c1", x"1e", x"26", x"40", x"a6", x"01", x"80", x"20", 
x"b1", x"ed", x"18", x"24", x"03", x"b7", x"ed", x"10", x"a6", x"02", x"80", x"20", x"b1", x"ed", x"17", x"24", 
x"03", x"b7", x"ed", x"11", x"20", x"59", x"81", x"7f", x"27", x"04", x"81", x"20", x"24", x"03", x"7e", x"fb", 
x"38", x"fe", x"ed", x"52", x"8d", x"17", x"b6", x"ed", x"10", x"4c", x"b1", x"ed", x"18", x"24", x"0d", x"b7", 
x"ed", x"10", x"fe", x"ed", x"52", x"08", x"ff", x"ed", x"52", x"7e", x"fa", x"fb", x"39", x"ff", x"ed", x"5d", 
x"37", x"b7", x"ed", x"5c", x"a7", x"00", x"b6", x"ed", x"5e", x"f6", x"ed", x"5d", x"b0", x"ed", x"16", x"f2", 
x"ed", x"15", x"f1", x"ed", x"13", x"26", x"03", x"b1", x"ed", x"14", x"25", x"0e", x"b7", x"ed", x"55", x"f7", 
x"ed", x"54", x"fe", x"ed", x"54", x"b6", x"ed", x"5c", x"a7", x"00", x"33", x"fe", x"ed", x"5d", x"39", x"b6", 
x"ed", x"18", x"4c", x"4c", x"b7", x"ed", x"5c", x"b6", x"ed", x"11", x"36", x"5f", x"37", x"b6", x"ed", x"10", 
x"5f", x"bb", x"ed", x"1a", x"f9", x"ed", x"19", x"b7", x"ed", x"53", x"f7", x"ed", x"52", x"74", x"ed", x"5c", 
x"24", x"0c", x"bb", x"ed", x"53", x"f9", x"ed", x"52", x"b7", x"ed", x"53", x"f7", x"ed", x"52", x"33", x"32", 
x"48", x"59", x"36", x"37", x"7d", x"ed", x"5c", x"26", x"e4", x"31", x"31", x"fe", x"ed", x"0e", x"bc", x"ed", 
x"0c", x"27", x"20", x"a6", x"00", x"fe", x"ed", x"22", x"81", x"fe", x"27", x"04", x"a1", x"01", x"26", x"07", 
x"3f", x"11", x"3f", x"04", x"fe", x"ed", x"22", x"81", x"fd", x"27", x"04", x"a1", x"00", x"26", x"04", x"3f", 
x"11", x"3f", x"11", x"b6", x"ed", x"53", x"f6", x"ed", x"52", x"8b", x"02", x"c9", x"00", x"36", x"17", x"c6", 
x"0e", x"8d", x"02", x"5c", x"32", x"7e", x"f4", x"7e", x"81", x"7f", x"26", x"0b", x"bd", x"fc", x"5b", x"fe", 
x"ed", x"52", x"86", x"20", x"7e", x"fa", x"8d", x"81", x"1e", x"26", x"04", x"c6", x"02", x"20", x"0a", x"81", 
x"1f", x"27", x"04", x"81", x"1b", x"26", x"0f", x"c6", x"01", x"ce", x"ed", x"59", x"a7", x"00", x"08", x"ff", 
x"ed", x"57", x"f7", x"ed", x"56", x"39", x"81", x"18", x"26", x"15", x"fe", x"ed", x"52", x"f6", x"ed", x"10", 
x"f1", x"ed", x"18", x"24", x"09", x"86", x"20", x"bd", x"fa", x"8d", x"08", x"5c", x"26", x"f2", x"39", x"81", 
x"0d", x"26", x"06", x"7f", x"ed", x"10", x"7e", x"fa", x"bf", x"81", x"0c", x"26", x"50", x"fe", x"ed", x"13", 
x"f6", x"ed", x"17", x"58", x"b6", x"ed", x"18", x"4c", x"4c", x"6f", x"00", x"08", x"4a", x"26", x"fa", x"5a", 
x"26", x"f2", x"8d", x"0f", x"7f", x"ed", x"10", x"7f", x"ed", x"11", x"fe", x"ed", x"19", x"ff", x"ed", x"52", 
x"7e", x"fa", x"fb", x"b6", x"ed", x"1a", x"f6", x"ed", x"19", x"bb", x"ed", x"16", x"f9", x"ed", x"15", x"b7", 
x"ed", x"21", x"f7", x"ed", x"20", x"fe", x"ed", x"20", x"0f", x"9f", x"0e", x"8e", x"bf", x"9f", x"c6", x"28", 
x"6f", x"00", x"32", x"32", x"a7", x"2a", x"08", x"5a", x"26", x"f6", x"9e", x"0e", x"39", x"81", x"0a", x"26", 
x"60", x"7f", x"ed", x"10", x"b6", x"ed", x"11", x"4c", x"b1", x"ed", x"17", x"24", x"06", x"b7", x"ed", x"11", 
x"7e", x"fa", x"bf", x"b6", x"ed", x"18", x"4c", x"4c", x"5f", x"bb", x"ed", x"1a", x"f9", x"ed", x"19", x"b7", 
x"ed", x"1a", x"f7", x"ed", x"19", x"b0", x"ed", x"16", x"f2", x"ed", x"15", x"f1", x"ed", x"13", x"26", x"03", 
x"b1", x"ed", x"14", x"24", x"ea", x"b6", x"ed", x"1a", x"f6", x"ed", x"19", x"bb", x"ed", x"16", x"f9", x"ed", 
x"15", x"b0", x"ed", x"18", x"c2", x"00", x"b7", x"ed", x"55", x"f7", x"ed", x"54", x"fe", x"ed", x"54", x"09", 
x"09", x"5f", x"bd", x"fb", x"70", x"bd", x"fb", x"b3", x"fe", x"ed", x"19", x"ff", x"ed", x"04", x"7e", x"fa", 
x"bf", x"81", x"09", x"26", x"12", x"b6", x"ed", x"10", x"8b", x"08", x"84", x"f8", x"b1", x"ed", x"18", x"24", 
x"03", x"b7", x"ed", x"10", x"7e", x"fa", x"bf", x"81", x"08", x"26", x"12", x"b6", x"ed", x"10", x"27", x"0a", 
x"7a", x"ed", x"10", x"fe", x"ed", x"52", x"09", x"ff", x"ed", x"52", x"7e", x"fa", x"fb", x"81", x"07", x"26", 
x"13", x"ce", x"00", x"c8", x"c6", x"64", x"5a", x"26", x"fd", x"b6", x"e6", x"2b", x"88", x"08", x"b7", x"e6", 
x"2b", x"09", x"26", x"f0", x"39", x"a6", x"00", x"27", x"05", x"3f", x"22", x"08", x"20", x"f7", x"39", x"5d", 
x"27", x"07", x"5a", x"27", x"3a", x"5a", x"27", x"1e", x"39", x"c6", x"0a", x"7d", x"e6", x"34", x"2a", x"0a", 
x"09", x"26", x"f8", x"5a", x"26", x"f5", x"86", x"01", x"20", x"26", x"b7", x"e6", x"35", x"86", x"34", x"b7", 
x"e6", x"36", x"86", x"3c", x"20", x"16", x"ce", x"00", x"00", x"ff", x"e6", x"36", x"ce", x"07", x"ff", x"ff", 
x"e6", x"34", x"86", x"34", x"b7", x"e6", x"37", x"86", x"3c", x"b7", x"e6", x"37", x"b7", x"e6", x"36", x"4f", 
x"ba", x"e6", x"34", x"7e", x"ff", x"f4", x"ce", x"00", x"08", x"5f", x"74", x"00", x"06", x"24", x"02", x"db", 
x"05", x"56", x"46", x"09", x"26", x"f4", x"7e", x"ff", x"f2", x"df", x"20", x"d7", x"22", x"97", x"23", x"26", 
x"07", x"5d", x"26", x"04", x"43", x"53", x"20", x"22", x"4f", x"5f", x"ce", x"00", x"11", x"49", x"59", x"90", 
x"23", x"d2", x"22", x"24", x"04", x"9b", x"23", x"d9", x"22", x"79", x"00", x"21", x"79", x"00", x"20", x"09", 
x"26", x"eb", x"73", x"00", x"21", x"73", x"00", x"20", x"de", x"20", x"7e", x"ff", x"f0", x"0f", x"c1", x"09", 
x"24", x"59", x"df", x"20", x"27", x"4f", x"30", x"df", x"22", x"b6", x"ee", x"1f", x"f6", x"ee", x"1e", x"90", 
x"21", x"d2", x"20", x"25", x"46", x"97", x"21", x"d7", x"20", x"d6", x"05", x"86", x"ff", x"5d", x"27", x"04", 
x"48", x"5a", x"20", x"f9", x"94", x"21", x"97", x"21", x"d6", x"20", x"b0", x"ee", x"1f", x"f2", x"ee", x"1e", 
x"9b", x"23", x"d9", x"22", x"24", x"25", x"97", x"23", x"d7", x"22", x"5a", x"f1", x"ee", x"1c", x"26", x"03", 
x"b1", x"ee", x"1d", x"25", x"16", x"de", x"22", x"32", x"a7", x"00", x"08", x"9c", x"20", x"26", x"f8", x"ff", 
x"ee", x"1e", x"de", x"22", x"35", x"fe", x"ee", x"1e", x"df", x"07", x"39", x"ce", x"00", x"00", x"df", x"07", 
x"39", x"0f", x"df", x"20", x"96", x"21", x"d6", x"20", x"f1", x"ee", x"1e", x"26", x"03", x"b1", x"ee", x"1f", 
x"23", x"2e", x"f1", x"ee", x"1a", x"26", x"03", x"b1", x"ee", x"1b", x"22", x"24", x"9f", x"22", x"35", x"fe", 
x"ee", x"1e", x"20", x"03", x"a6", x"00", x"36", x"09", x"9c", x"22", x"26", x"f8", x"96", x"21", x"d6", x"20", 
x"b0", x"ee", x"1f", x"f2", x"ee", x"1e", x"97", x"08", x"d7", x"07", x"de", x"20", x"ff", x"ee", x"1e", x"39", 
x"ce", x"00", x"00", x"df", x"07", x"39", x"fe", x"ee", x"1e", x"ff", x"ee", x"1a", x"39", x"0f", x"ee", x"00", 
x"df", x"22", x"09", x"df", x"20", x"de", x"07", x"ee", x"02", x"df", x"26", x"97", x"08", x"d7", x"07", x"4d", 
x"26", x"03", x"5d", x"27", x"45", x"9b", x"21", x"d9", x"20", x"97", x"21", x"d7", x"20", x"9f", x"0e", x"96", 
x"21", x"d6", x"20", x"90", x"23", x"d2", x"22", x"9b", x"27", x"d9", x"26", x"97", x"25", x"d7", x"24", x"96", 
x"26", x"91", x"22", x"26", x"04", x"96", x"27", x"91", x"23", x"23", x"0f", x"9e", x"24", x"de", x"20", x"08", 
x"09", x"a6", x"00", x"36", x"9c", x"22", x"26", x"f8", x"20", x"0e", x"9e", x"22", x"de", x"26", x"34", x"09", 
x"08", x"32", x"a7", x"00", x"9c", x"24", x"26", x"f8", x"9e", x"0e", x"39", x"0f", x"16", x"54", x"d7", x"0d", 
x"c6", x"ed", x"d7", x"0c", x"de", x"0c", x"e6", x"80", x"25", x"04", x"54", x"54", x"54", x"54", x"c4", x"0f", 
x"d7", x"05", x"c6", x"77", x"48", x"59", x"97", x"0d", x"d7", x"0c", x"de", x"0c", x"ee", x"00", x"df", x"07", 
x"39", x"0f", x"9f", x"0e", x"35", x"31", x"97", x"0a", x"44", x"97", x"0d", x"86", x"ed", x"97", x"0c", x"de", 
x"0c", x"86", x"0f", x"24", x"02", x"86", x"f0", x"a4", x"80", x"97", x"0b", x"17", x"84", x"0f", x"25", x"04", 
x"48", x"48", x"48", x"48", x"9a", x"0b", x"a7", x"80", x"86", x"77", x"d6", x"0a", x"58", x"49", x"d7", x"0d", 
x"97", x"0c", x"de", x"0c", x"af", x"00", x"9e", x"0e", x"39", x"0f", x"fe", x"ee", x"1c", x"df", x"07", x"9f", 
x"0e", x"7a", x"00", x"0e", x"bb", x"ee", x"1d", x"f9", x"ee", x"1c", x"d1", x"0e", x"26", x"02", x"91", x"0f", 
x"24", x"07", x"f7", x"ee", x"1c", x"b7", x"ee", x"1d", x"39", x"7f", x"00", x"05", x"7f", x"00", x"06", x"39", 
x"0f", x"fe", x"ee", x"1c", x"9f", x"0e", x"96", x"0f", x"d6", x"0e", x"5a", x"b0", x"ee", x"1d", x"f2", x"ee", 
x"1c", x"24", x"02", x"5f", x"4f", x"7e", x"ff", x"f0", x"0f", x"8c", x"00", x"00", x"26", x"06", x"ce", x"ff", 
x"f6", x"df", x"07", x"5f", x"30", x"e7", x"02", x"d6", x"07", x"96", x"08", x"e7", x"08", x"a7", x"09", x"a6", 
x"03", x"97", x"04", x"e6", x"04", x"a6", x"05", x"ee", x"06", x"7e", x"ff", x"f0", x"f2", x"0b", x"f2", x"0b", 
x"00", x"00", x"00", x"00", x"00", x"00", x"f2", x"18", x"00", x"00", x"00", x"00", x"00", x"00", x"f2", x"ab", 
x"00", x"00", x"00", x"00", x"00", x"00", x"be", x"00", x"01", x"00", x"be", x"00", x"f3", x"72", x"f3", x"82", 
x"f3", x"c5", x"f4", x"85", x"f4", x"99", x"f4", x"a6", x"f4", x"ba", x"f4", x"bf", x"f9", x"4a", x"f9", x"5a", 
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"f9", x"86", x"f9", x"c6", 
x"fa", x"16", x"fc", x"85", x"00", x"00", x"00", x"00", x"fc", x"8f", x"00", x"00", x"fc", x"d6", x"fc", x"e9", 
x"fd", x"1d", x"fd", x"81", x"fd", x"c6", x"fd", x"cd", x"fe", x"2b", x"fe", x"51", x"00", x"00", x"00", x"00", 
x"00", x"00", x"00", x"00", x"00", x"00", x"fe", x"89", x"fe", x"b0", x"fe", x"c8", x"6f", x"03", x"02", x"09", 
x"2a", x"ff", x"50", x"ff", x"80", x"00", x"00", x"00", x"01", x"01", x"00", x"13", x"03", x"06", x"07", x"00", 
x"07", x"20", x"07", x"3f", x"28", x"30", x"05", x"26", x"00", x"19", x"1f", x"00", x"07", x"20", x"07", x"f0", 
x"00", x"f0", x"00", x"04", x"1a", x"00", x"3e", x"24", x"38", x"00", x"7e", x"08", x"80", x"0a", x"28", x"43", 
x"29", x"20", x"53", x"6f", x"66", x"74", x"77", x"61", x"72", x"65", x"20", x"52", x"44", x"4c", x"20", x"31", 
x"39", x"38", x"37", x"2d", x"38", x"39", x"2c", x"20", x"49", x"76", x"6f", x"20", x"4e", x"65", x"6e", x"6f", 
x"76", x"0a", x"20", x"26", x"20", x"4f", x"72", x"6c", x"69", x"6e", x"20", x"53", x"68", x"6f", x"70", x"6f", 
x"76", x"20", x"2d", x"20", x"45", x"61", x"67", x"6c", x"65", x"20", x"73", x"6f", x"66", x"74", x"77", x"61", 
x"72", x"65", x"0a", x"00", x"ff", x"ff", x"ff", x"89", x"07", x"1e", x"30", x"20", x"8f", x"ba", x"ab", x"a4", 
x"a8", x"ad", x"20", x"36", x"30", x"31", x"20", x"00", x"b4", x"61", x"00", x"00", x"b4", x"61", x"02", x"32", 
x"df", x"07", x"d7", x"05", x"97", x"06", x"39", x"00", x"f1", x"53", x"f1", x"89", x"f1", x"47", x"f0", x"06" 
);
begin
	data <= rom_data(conv_integer(addr));
end basic;
