--===========================================================================--
--
--  S Y N T H E Z I A B L E    SWTBUG ROM   C O R E
--
--  www.OpenCores.Org - December 2002
--  This core adheres to the GNU public license  
--
-- File name      : swtbug.vhd
--
-- entity name    : rombios_rom
--
-- Purpose        : Implements a 1K x 8 ROM containing the
--                  SWTBUG rombios program for the SWTPC 6800
--                  
-- Dependencies   : ieee.Std_Logic_1164
--                  ieee.std_logic_unsigned
--                  ieee.std_logic_arith
--
-- Author         : John E. Kent      
--
--===========================================================================----
--
-- Revision History:
--
-- Date:          Revision         Author
-- 22 Sep 2002    0.1              John Kent
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity rombios_rom is
  port (
    cs     : in  std_logic;
    addr   : in  std_logic_vector(9 downto 0);
    data   : out std_logic_vector(7 downto 0)
  );
end;

architecture basic of rombios_rom is
  constant width   : integer := 8;
  constant memsize : integer := 4096;

  type rom_array is array(0 to memsize-1) of std_logic_vector(width-1 downto 0);

  constant rom_data : rom_array :=
(
"11111110",
"10100000",
"00000000",
"01101110",
"00000000",
"10001101",
"01000000",
"01101110",
"00000000",
"00010000",
"00010110",
"00000100",
"10111101",
"11100011",
"00110100",
"10001101",
"01100111",
"10000001",
"01010011",
"00100110",
"11111010",
"10001101",
"01100001",
"10000001",
"00111001",
"00100111",
"00101001",
"10000001",
"00110001",
"00100110",
"11110000",
"01111111",
"10100000",
"00001111",
"10001101",
"00110001",
"10000000",
"00000010",
"10110111",
"10100000",
"01000111",
"10001101",
"00011100",
"10001101",
"00101000",
"01111010",
"10100000",
"01000111",
"00100111",
"00001001",
"10100111",
"00000000",
"10100001",
"00000000",
"00100110",
"00001000",
"00001000",
"00100000",
"11110000",
"01111100",
"10100000",
"00001111",
"00100111",
"11001111",
"10000110",
"00111111",
"10001101",
"00110001",
"01111110",
"11100010",
"11010100",
"10001101",
"00001100",
"10110111",
"10100000",
"00001101",
"10001101",
"00000111",
"10110111",
"10100000",
"00001110",
"11111110",
"10100000",
"00001101",
"00111001",
"10001101",
"01010011",
"01001000",
"01001000",
"01001000",
"01001000",
"00010110",
"10001101",
"01001100",
"00011011",
"00010110",
"11111011",
"10100000",
"00001111",
"11110111",
"10100000",
"00001111",
"00111001",
"01000100",
"01000100",
"01000100",
"01000100",
"10000100",
"00001111",
"10001011",
"00110000",
"10000001",
"00111001",
"00100011",
"00000010",
"10001011",
"00000111",
"01111110",
"11100001",
"11010001",
"01111110",
"11100001",
"10101100",
"10001101",
"11111000",
"00001000",
"10100110",
"00000000",
"10000001",
"00000100",
"00100110",
"11110111",
"00111001",
"01111110",
"11100001",
"01001010",
"10001101",
"10111101",
"11001110",
"11100001",
"10011101",
"10001101",
"11101111",
"11001110",
"10100000",
"00001101",
"10001101",
"00110100",
"11111110",
"10100000",
"00001101",
"10001101",
"00110001",
"10001101",
"00110001",
"10001101",
"11011011",
"10000001",
"00100000",
"00100111",
"11111010",
"10000001",
"00001101",
"00100111",
"11100000",
"10000001",
"01011110",
"00100000",
"00101100",
"00000001",
"10001101",
"11001100",
"10000000",
"00110000",
"00101011",
"01001100",
"10000001",
"00001001",
"00101111",
"00001010",
"10000001",
"00010001",
"00101011",
"01000100",
"10000001",
"00010110",
"00101110",
"01000000",
"10000000",
"00000111",
"00111001",
"10100110",
"00000000",
"10001101",
"10100100",
"10100110",
"00000000",
"00001000",
"00100000",
"10100011",
"10001101",
"11110101",
"10001101",
"11110011",
"10000110",
"00100000",
"00100000",
"10100101",
"10001110",
"10100000",
"01000010",
"00100000",
"00101100",
"00100110",
"00000111",
"00001001",
"00001001",
"11111111",
"10100000",
"00001101",
"00100000",
"10101100",
"11111111",
"10100000",
"00001101",
"00100000",
"00000010",
"00100000",
"01101101",
"10000001",
"00110000",
"00100101",
"10100001",
"10000001",
"01000110",
"00100010",
"10011101",
"10001101",
"10111101",
"10111101",
"11100000",
"01010111",
"00001001",
"10100111",
"00000000",
"10100001",
"00000000",
"00100111",
"10010001",
"01111110",
"11100000",
"01000000",
"10111110",
"10100000",
"00001000",
"00100000",
"01001001",
"10111111",
"10100000",
"00001000",
"10000110",
"11111111",
"10111101",
"11100011",
"00001000",
"11001110",
"10000000",
"00000100",
"10111101",
"11100010",
"10000100",
"10100110",
"00000000",
"10100001",
"00000010",
"00100000",
"00000010",
"00100000",
"00011001",
"00100110",
"00111001",
"10000110",
"00000011",
"10100111",
"00000000",
"10000110",
"00010001",
"10100111",
"00000000",
"00100000",
"00101111",
"00000001",
"10111111",
"10100000",
"00001000",
"00110000",
"01101101",
"00000110",
"00100110",
"00000010",
"01101010",
"00000101",
"01101010",
"00000110",
"11001110",
"11100001",
"10011101",
"10111101",
"11100000",
"01111110",
"11111110",
"10100000",
"00001000",
"00001000",
"10001101",
"10001110",
"10001101",
"10001100",
"10001101",
"10001010",
"10001101",
"10000110",
"10001101",
"10000100",
"11001110",
"10100000",
"00001000",
"10111101",
"11100000",
"11001000",
"11111110",
"10100000",
"00010010",
"10001100",
"11100001",
"00100011",
"00100111",
"00011001",
"10001110",
"10100000",
"01000010",
"11001110",
"10000000",
"00000100",
"11111111",
"10100000",
"00001010",
"01111111",
"10100000",
"00001100",
"10001101",
"01110011",
"00100111",
"00000011",
"10111101",
"11100010",
"01111101",
"10111101",
"11100011",
"01010011",
"10111101",
"11100011",
"01000111",
"11001110",
"11100001",
"10011100",
"10111101",
"11100000",
"01111110",
"10001101",
"00111001",
"11001110",
"11100011",
"11010001",
"10100001",
"00000000",
"00100110",
"00000111",
"10111101",
"11100000",
"11001100",
"11101110",
"00000001",
"01101110",
"00000000",
"00001000",
"00001000",
"00001000",
"10001100",
"11100011",
"11111000",
"00100110",
"11101101",
"00100000",
"10111111",
"11111110",
"10100000",
"00010010",
"01101110",
"00000000",
"01010011",
"00111001",
"00000100",
"00001101",
"00001010",
"00010101",
"00000000",
"00000000",
"00000000",
"01010011",
"00110001",
"00000100",
"00010011",
"00001101",
"00001010",
"00010101",
"00000000",
"00000000",
"00000000",
"00100100",
"00000100",
"00100000",
"01001100",
"11111110",
"10100000",
"00000110",
"01101110",
"00000000",
"00100000",
"01000000",
"10111101",
"11100000",
"01000111",
"11111111",
"10100000",
"00000100",
"10111101",
"11100000",
"01000111",
"10111101",
"11100000",
"01010101",
"00010110",
"10100110",
"00000000",
"11111111",
"10100000",
"00001101",
"00010001",
"00100111",
"00000010",
"00100000",
"00100001",
"11001110",
"11100001",
"10011101",
"10111101",
"11100000",
"01111110",
"11001110",
"10100000",
"00001101",
"00100000",
"00010000",
"00111011",
"00100000",
"00111010",
"11111111",
"10100000",
"00010000",
"11111110",
"10100000",
"00001010",
"00110111",
"11100110",
"00000001",
"11100001",
"00000011",
"00110011",
"00111001",
"10111101",
"11100000",
"11001000",
"11111110",
"10100000",
"00001101",
"10111100",
"10100000",
"00000100",
"00100111",
"10011110",
"00001000",
"00100000",
"11001101",
"10001101",
"00000110",
"10000100",
"01111111",
"00111001",
"00110001",
"00110001",
"00110001",
"00110111",
"10001101",
"11011010",
"00100110",
"00101000",
"10000110",
"00010101",
"10100111",
"00000000",
"10100110",
"00000000",
"01000111",
"00100100",
"11111011",
"10100110",
"00000001",
"11110110",
"10100000",
"00001100",
"00100111",
"00000111",
"00100000",
"00010001",
"00110111",
"10001101",
"11000011",
"00100110",
"00101110",
"11000110",
"00010001",
"11100111",
"00000000",
"11100110",
"00000000",
"01010111",
"01010111",
"00100100",
"11111010",
"10100111",
"00000001",
"00110011",
"11111110",
"10100000",
"00010000",
"00111001",
"10100110",
"00000000",
"00101011",
"11111100",
"10001101",
"00111010",
"11000110",
"00000100",
"11100111",
"00000010",
"01011000",
"10001101",
"00101010",
"00001101",
"01101001",
"00000000",
"01000110",
"01011010",
"00100110",
"11110111",
"10001101",
"00100001",
"11110110",
"10100000",
"00001100",
"00100111",
"00010011",
"00100000",
"11011110",
"10001101",
"00100011",
"11000110",
"00001010",
"01101010",
"00000000",
"10001101",
"00010110",
"10001101",
"00010000",
"10100111",
"00000000",
"00001101",
"01000110",
"01011010",
"00100110",
"11110111",
"11100110",
"00000010",
"01011000",
"00101010",
"11001000",
"10001101",
"00000010",
"00100000",
"11000100",
"01101101",
"00000010",
"00101010",
"11111100",
"01101100",
"00000010",
"01101010",
"00000010",
"00111001",
"01101111",
"00000010",
"10001101",
"11110111",
"00100000",
"11110001",
"10001101",
"10000011",
"00010110",
"01111111",
"10100000",
"00001011",
"11111110",
"10100000",
"00001010",
"10001101",
"00010000",
"10001101",
"00000111",
"11001110",
"11100011",
"11101111",
"00010111",
"01111110",
"11100001",
"01110110",
"10000110",
"00110100",
"10100111",
"00000011",
"10100111",
"00000010",
"00111001",
"01101100",
"00000000",
"10000110",
"00000111",
"10100111",
"00000001",
"01101100",
"00000000",
"10100111",
"00000010",
"00111001",
"01111111",
"10000000",
"00010100",
"10001101",
"00101110",
"11000110",
"00001011",
"10001101",
"00100101",
"11100110",
"00000100",
"11000101",
"00000001",
"00100110",
"11111010",
"01101111",
"00000110",
"10001101",
"00011101",
"11000110",
"10011100",
"10001101",
"00010111",
"11001110",
"00100100",
"00000000",
"11000101",
"00000010",
"00100111",
"00000110",
"10110110",
"10000000",
"00011011",
"10100111",
"00000000",
"00001000",
"11110110",
"10000000",
"00011000",
"11000101",
"00000001",
"00100110",
"11101111",
"01111110",
"00100100",
"00000000",
"11100111",
"00000100",
"10001101",
"00000000",
"00111001",
"11001110",
"11111111",
"11111111",
"00001001",
"10001100",
"10000000",
"00010100",
"00100110",
"11111010",
"00111001",
"11001110",
"11100000",
"00001001",
"10111101",
"11100000",
"01111110",
"10001101",
"11110001",
"10111101",
"11100011",
"01000111",
"00100000",
"01011000",
"11001110",
"11100001",
"00100011",
"10111100",
"10100000",
"00010010",
"00100111",
"00011010",
"00001000",
"10001101",
"00110010",
"10111101",
"11100000",
"01000111",
"11111111",
"10100000",
"00010100",
"10100110",
"00000000",
"10110111",
"10100000",
"00010110",
"10000110",
"00111111",
"10100111",
"00000000",
"11001110",
"11100001",
"00100011",
"10001101",
"00011110",
"01111110",
"11100001",
"01101011",
"11111110",
"10100000",
"00010100",
"10110110",
"10100000",
"00010110",
"10100111",
"00000000",
"11001110",
"11100001",
"00100100",
"00100000",
"11011010",
"10110111",
"10100000",
"01000011",
"11111110",
"10100000",
"00010010",
"10001100",
"11100001",
"00100011",
"00100111",
"00000110",
"11001110",
"11100001",
"00100100",
"11111111",
"10100000",
"00010010",
"00111001",
"10001101",
"01011010",
"00100000",
"00001111",
"11001110",
"10100000",
"01001001",
"11111111",
"10100000",
"00000100",
"00001001",
"10001101",
"01010010",
"11001110",
"11100001",
"10010000",
"10111101",
"11100000",
"01111110",
"10001101",
"00100100",
"10001101",
"10010001",
"01111110",
"11100001",
"01010010",
"01110011",
"10100000",
"00001100",
"10000110",
"00010001",
"11000110",
"00100000",
"10001101",
"00011010",
"10111101",
"11100001",
"11011001",
"00100111",
"00000100",
"10000110",
"00111100",
"10100111",
"00000011",
"00111001",
"10000110",
"00010011",
"11000110",
"00010000",
"00100000",
"00001010",
"10000110",
"00010010",
"11000110",
"00000100",
"00100000",
"00000100",
"10000110",
"00010100",
"11000110",
"00001000",
"10111101",
"11100000",
"01110101",
"10111101",
"11100001",
"11010110",
"00100111",
"00010110",
"10000110",
"00000010",
"11001010",
"00000001",
"10001101",
"00001100",
"10001101",
"00001000",
"10000110",
"00000010",
"11000110",
"00000001",
"11100111",
"00000000",
"10001101",
"00000010",
"10000110",
"00000110",
"10100111",
"00000001",
"11100111",
"00000000",
"00111001",
"11111110",
"10100000",
"00000010",
"11111111",
"10100000",
"01000100",
"10001101",
"11001111",
"10110110",
"10100000",
"00000101",
"10110000",
"10100000",
"01000101",
"11110110",
"10100000",
"00000100",
"11110010",
"10100000",
"01000100",
"00100110",
"00000100",
"10000001",
"00010000",
"00100101",
"00000010",
"10000110",
"00001111",
"10001011",
"00000100",
"10110111",
"10100000",
"01000111",
"10000000",
"00000011",
"10110111",
"10100000",
"01000110",
"11001110",
"11100001",
"10010011",
"10111101",
"11100000",
"01111110",
"01011111",
"11001110",
"10100000",
"01000111",
"10001101",
"00100100",
"11001110",
"10100000",
"01000100",
"10001101",
"00011111",
"10001101",
"00011101",
"11111110",
"10100000",
"01000100",
"10001101",
"00011000",
"01111010",
"10100000",
"01000110",
"00100110",
"11111001",
"11111111",
"10100000",
"01000100",
"01010011",
"00110111",
"00110000",
"10001101",
"00001011",
"00110011",
"11111110",
"10100000",
"01000100",
"00001001",
"10111100",
"10100000",
"00000100",
"00100110",
"10110011",
"00111001",
"11101011",
"00000000",
"01111110",
"11100000",
"10111111",
"01000111",
"11100001",
"11010000",
"01011010",
"11000000",
"00000000",
"01001101",
"11100000",
"10001000",
"01000110",
"11100001",
"10101110",
"01010010",
"11100001",
"00110000",
"01001010",
"11100000",
"00000101",
"01000011",
"11100010",
"11001100",
"01000100",
"11100010",
"10001111",
"01000010",
"11100010",
"11011001",
"01001111",
"11100010",
"01101001",
"01010000",
"11100011",
"00011010",
"01001100",
"11100000",
"00001100",
"01000101",
"11100011",
"00011110",
"11100000",
"00000000",
"11100001",
"10001011",
"11100001",
"10100111",
"11100000",
"11010000"
);
begin
   data <= rom_data(conv_integer(addr));
end;

